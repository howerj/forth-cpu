-- SPI, AD5641 Interface
library ieee,work,std;
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;

entity spi_ad5641 is
  port(

      );
end entity;

architecture rtl of spi_ad5641 is

begin


end architecture;
