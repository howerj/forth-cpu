../../../vhd/gptimer.vhd