-- SPI, AD5641 Interface
