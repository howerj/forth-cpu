spi_ad5641/spi_ad5641.vhd