-- Richard James Howe.
--  I/O control module
--
-- @author     Richard James Howe.
-- @copyright    Copyright 2013 Richard James Howe.
-- @license    LGPL    
-- @email      howe.r.j.89@gmail.com
library ieee,work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity io is
  port(
      clk:  in std_logic := 'X'
      );
end;

architecture behav of io is
begin


end architecture;
