../../../vhdl/uart.vhd