../../../vhdl/gptimer.vhd