spi_ad5641/shift_reg_16.vhd