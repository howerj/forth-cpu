-- Timer
